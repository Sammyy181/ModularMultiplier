`timescale 1ns / 1ps

module rectKaratsuba(
    input wire clock,
    input wire in_valid,
    input wire [255:0] X,
    input wire [255:0] Y,
    input wire reset,
    output reg [511:0] P,
    output reg out_valid,
    output reg [41:0] Z0_S1, Z3_S1, Z4_S1, Z6_S1, Z7_S1, Z8_S1, Z9_S1,
                Z10_S1, Z11_S1, Z13_S1, Z14_S1,  Z17_S1,
                Z20_S1, Z23_S1, Z24_S1, Z25_S1, Z26_S1, Z27_S1, Z28_S1,
                Z30_S1, Z31_S1, Z32_S1, Z33_S1, Z34_S1, Z35_S1, Z37_S1, Z38_S1,
                Z41_S1, Z44_S1, Z45_S1, Z47_S1, Z48_S1, Z49_S1,
                Z50_S1, Z51_S1, Z52_S1, Z54_S1, Z55_S1, Z56_S1, Z57_S1, Z58_S1, Z59_S1,
                Z62_S1, Z65_S1, Z68_S1, Z69_S1,
                Z71_S1, Z72_S1, Z75_S1,
    output reg [33:0] Z73_S1, Z76_S1, Z79_S1,
    output reg [27:0] Z74_S1, Z78_S1,
    output reg [19:0] Z82_S1
    );

    // 1st Cycle
    /*
    reg [41:0] Z0_S1, Z3_S1, Z4_S1, Z6_S1, Z7_S1, Z8_S1, Z9_S1,
                Z10_S1, Z11_S1, Z13_S1, Z14_S1,  Z17_S1,
                Z20_S1, Z23_S1, Z24_S1, Z25_S1, Z26_S1, Z27_S1, Z28_S1,
                Z30_S1, Z31_S1, Z32_S1, Z33_S1, Z34_S1, Z35_S1, Z37_S1, Z38_S1,
                Z41_S1, Z44_S1, Z45_S1, Z47_S1, Z48_S1, Z49_S1,
                Z50_S1, Z51_S1, Z52_S1, Z54_S1, Z55_S1, Z56_S1, Z57_S1, Z58_S1, Z59_S1,
                Z62_S1, Z65_S1, Z68_S1, Z69_S1,
                Z71_S1, Z72_S1, Z75_S1;
    reg [33:0] Z73_S1, Z76_S1, Z79_S1;
    reg [27:0] Z74_S1, Z78_S1;
    reg [19:0] Z82_S1;
    */
    reg S1_valid;

    always @(posedge clock) begin
        if(reset) begin
            P <= 512'b0;
            S1_valid <= 1'b0;
            out_valid <= 1'b0;
        end

        // 1st Cycle
        Z0_S1[41:0] <= X[17:0] * Y[23:0];
        Z3_S1[41:0] <= X[35:18] * Y[23:0];
        Z4_S1[41:0] <= X[17:0] * Y[47:24];
        Z6_S1[41:0] <= X[53:36] * Y[23:0];
        Z7_S1[41:0] <= X[35:18] * Y[47:24];
        Z8_S1[41:0] <= X[17:0] * Y[71:48];
        Z9_S1[41:0] <= X[71:54] * Y[23:0];
        Z10_S1[41:0] <= X[53:36] * Y[47:24];
        Z11_S1[41:0] <= X[35:18] * Y[71:48];
        Z13_S1[41:0] <= X[71:54] * Y[47:24];
        Z14_S1[41:0] <= X[53:36] * Y[71:48];
        Z17_S1[41:0] <= X[71:54] * Y[71:48];
        Z20_S1[41:0] <= X[89:72] * Y[71:48];
        Z23_S1[41:0] <= X[107:90] * Y[71:48];
        Z24_S1[41:0] <= X[89:72] * Y[95:72];
        Z25_S1[41:0] <= X[71:54] * Y[119:96];
        Z26_S1[41:0] <= X[125:108] * Y[71:48];
        Z27_S1[41:0] <= X[107:90] * Y[95:72];
        Z28_S1[41:0] <= X[89:72] * Y[95:72];
        Z30_S1[41:0] <= X[125:108] * Y[95:72];
        Z31_S1[41:0] <= X[107:90] * Y[119:96];
        Z32_S1[41:0] <= X[89:72] * Y[143:120];
        Z33_S1[41:0] <= X[143:126] * Y[95:72];
        Z34_S1[41:0] <= X[125:108] * Y[119:96];
        Z35_S1[41:0] <= X[107:90] * Y[143:120];
        Z37_S1[41:0] <= X[143:126] * Y[119:96];
        Z38_S1[41:0] <= X[125:108] * Y[143:120];
        Z41_S1[41:0] <= X[143:126] * Y[143:120];
        Z44_S1[41:0] <= X[161:144] * Y[143:120];
        Z45_S1[41:0] <= X[143:126] * Y[167:144];
        Z47_S1[41:0] <= X[179:162] * Y[143:120];
        Z48_S1[41:0] <= X[161:144] * Y[167:144];
        Z49_S1[41:0] <= X[179:162] * Y[191:168];
        Z50_S1[41:0] <= X[197:180] * Y[143:120];
        Z51_S1[41:0] <= X[179:162] * Y[167:144];
        Z52_S1[41:0] <= X[161:144] * Y[191:168];
        Z54_S1[41:0] <= X[197:180] * Y[167:144];
        Z55_S1[41:0] <= X[179:162] * Y[191:168];
        Z56_S1[41:0] <= X[161:144] * Y[215:192];
        Z57_S1[41:0] <= X[215:198] * Y[167:144];
        Z58_S1[41:0] <= X[197:180] * Y[191:168];
        Z59_S1[41:0] <= X[179:162] * Y[215:192];
        Z62_S1[41:0] <= X[197:180] * Y[215:192];
        Z65_S1[41:0] <= X[215:198] * Y[215:192];
        Z68_S1[41:0] <= X[233:216] * Y[215:192];
        Z69_S1[41:0] <= X[215:198] * Y[239:216];
        Z71_S1[41:0] <= X[251:234] * Y[215:192];
        Z72_S1[41:0] <= X[233:216] * Y[239:216];
        Z73_S1[33:0] <= X[215:198] * Y[255:240];
        Z74_S1[27:0] <= X[255:252] * Y[215:192];
        Z75_S1[41:0] <= X[251:234] * Y[239:216];
        Z76_S1[33:0] <= X[233:216] * Y[255:240];
        Z78_S1[27:0] <= X[255:252] * Y[239:216];
        Z79_S1[33:0] <= X[251:234] * Y[255:240];
        Z82_S1[19:0] <= X[255:252] * Y[255:240];
        S1_valid <= in_valid;
    end

endmodule