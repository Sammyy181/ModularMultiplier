`timescale 1ns/1ps

module fastKaratsuba(
    input wire clock,
    input wire reset,
    input wire [255:0] X,
    input wire [255:0] Y,
    input wire in_valid,
    output reg [511:0] P,
    output reg out_valid,
    output reg [39:0] Z0_S1, Z2_S1, Z3_S1, Z4_S1, Z5_S1, Z7_S1, Z8_S1, Z9_S1,
                Z10_S1, Z12_S1, Z14_S1, Z15_S1, Z16_S1, Z17_S1, Z19_S1,
                Z20_S1, Z21_S1, Z22_S1, Z24_S1, Z26_S1, Z27_S1, Z28_S1, Z29_S1,
                Z31_S1, Z32_S1, Z33_S1, Z34_S1, Z36_S1, Z38_S1, Z39_S1,
                Z40_S1, Z41_S1, Z43_S1, Z44_S1, Z45_S1, Z46_S1, Z48_S1,
                Z50_S1, Z51_S1, Z52_S1, Z53_S1, Z55_S1, Z57_S1,
    output reg [31:0] Z56_S1, Z58_S1, Z60_S1,
    output reg [42:0] M6_S1, M8_S1, M9_S1, M10_S1, M11_S1, M12_S1, M13_S1, M14_S1, M15_S1, M16_S1, M17_S1, M18_0S1, M18_1S1, M19_S1,
                M20_0S1, M20_1S1, M21_0S1, M21_1S1, M22_0S1, M22_1S1, M23_0S1, M23_1S1, M24_0S1, M24_1S1, M25_0S1, M25_1S1,
                M26_0S1, M26_1S1, M27_0S1, M27_1S1, M28_0S1, M28_1S1, M29_0S1, M29_1S1, M30_0S1, M30_1S1, M30_2S1, M31_0S1,
                M31_1S1, M32_0S1, M32_1S1, M33_0S1, M33_1S1, M34_0S1, M34_1S1, M35_0S1, M35_1S1, M36_0S1, M36_1S1, M37_0S1,
                M37_1S1, M38_0S1, M38_1S1, M39_0S1, M39_1S1, M40_0S1, M40_1S1, M41_S1, M42_0S1, M42_1S1, M43_S1, M44_S1, M45_S1,
                M46_S1, M47_S1, M48_S1, M49_S1, M50_S1, M51_S1, M52_S1, M54_S1
);

    // Cycle 1
    /*
    reg [39:0] Z0_S1, Z2_S1, Z3_S1, Z4_S1, Z5_S1, Z7_S1, Z8_S1, Z9_S1,
                Z10_S1, Z12_S1, Z14_S1, Z15_S1, Z16_S1, Z17_S1, Z19_S1,
                Z20_S1, Z21_S1, Z22_S1, Z24_S1, Z26_S1, Z27_S1, Z28_S1, Z29_S1,
                Z31_S1, Z32_S1, Z33_S1, Z34_S1, Z36_S1, Z38_S1, Z39_S1,
                Z40_S1, Z41_S1, Z43_S1, Z44_S1, Z45_S1, Z46_S1, Z48_S1,
                Z50_S1, Z51_S1, Z52_S1, Z53_S1, Z55_S1, Z57_S1;
    reg [31:0] Z56_S1, Z58_S1, Z60_S1;

    reg [42:0] M6_S1, M8_S1, M9_S1, M10_S1, M11_S1, M12_S1, M13_S1, M14_S1, M15_S1, M16_S1, M17_S1, M18_0S1, M18_1S1, M19_S1,
                M20_0S1, M20_1S1, M21_0S1, M21_1S1, M22_0S1, M22_1S1, M23_0S1, M23_1S1, M24_0S1, M24_1S1, M25_0S1, M25_1S1,
                M26_0S1, M26_1S1, M27_0S1, M27_1S1, M28_0S1, M28_1S1, M29_0S1, M29_1S1, M30_0S1, M30_1S1, M30_2S1, M31_0S1,
                M31_1S1, M32_0S1, M32_1S1, M33_0S1, M33_1S1, M34_0S1, M34_1S1, M35_0S1, M35_1S1, M36_0S1, M36_1S1, M37_0S1,
                M37_1S1, M38_0S1, M38_1S1, M39_0S1, M39_1S1, M40_0S1, M40_1S1, M41_S1, M42_0S1, M42_1S1, M43_S1, M44_S1, M45_S1,
                M46_S1, M47_S1, M48_S1, M49_S1, M50_S1, M51_S1, M52_S1, M54_S1; 
    */
    reg S1_valid;

    // Cycle 2
    reg S2_valid;

    always @(posedge clock) begin
        if(reset) begin
            P <= 256'b0;
            S1_valid <= 1'b0;
            out_valid <= 1'b0;
        end
        else begin

            // Cycle 1
            Z0_S1 <= X[15:0] * Y[23:0];
            Z2_S1 <= X[31:16] * Y[23:0];
            Z3_S1 <= X[15:0] * Y[47:24];
            Z4_S1 <= X[47:32] * Y[23:0];
            Z5_S1 <= X[31:16] * Y[47:24];
            Z7_S1 <= X[47:32] * Y[47:24];
            Z8_S1 <= X[31:16] * Y[71:48];
            Z9_S1 <= X[63:48] * Y[47:24];
            Z10_S1 <= X[47:32] * Y[71:48];
            Z12_S1 <= X[63:48] * Y[71:48];
            Z14_S1 <= X[79:64] * Y[71:48];
            Z15_S1 <= X[63:48] * Y[95:72];
            Z16_S1 <= X[97:80] * Y[71:48];
            Z17_S1 <= X[79:64] * Y[95:72];
            Z19_S1 <= X[95:80] * Y[95:72];
            Z20_S1 <= X[79:64] * Y[119:96];
            Z21_S1 <= X[111:96] * Y[95:72];
            Z22_S1 <= X[95:80] * Y[119:96];
            Z24_S1 <= X[111:96] * Y[119:96];
            Z26_S1 <= X[127:112] * Y[119:96];
            Z27_S1 <= X[111:96] * Y[143:120];
            Z28_S1 <= X[143:128] * Y[119:96];
            Z29_S1 <= X[127:112] * Y[143:120];
            Z31_S1 <= X[143:128] * Y[143:120];
            Z32_S1 <= X[127:112] * Y[167:144];
            Z33_S1 <= X[159:144] * Y[143:120];
            Z34_S1 <= X[143:128] * Y[167:144];
            Z36_S1 <= X[159:144] * Y[167:144];
            Z38_S1 <= X[175:160] * Y[167:144];
            Z39_S1 <= X[159:144] * Y[191:168];
            Z40_S1 <= X[191:176] * Y[167:144];
            Z41_S1 <= X[175:160] * Y[191:168];
            Z43_S1 <= X[191:176] * Y[191:168];
            Z44_S1 <= X[175:160] * Y[215:192];
            Z45_S1 <= X[207:192] * Y[191:168];
            Z46_S1 <= X[191:176] * Y[215:192];
            Z48_S1 <= X[207:192] * Y[215:192];
            Z50_S1 <= X[223:208] * Y[215:192];
            Z51_S1 <= X[207:192] * Y[239:216];
            Z52_S1 <= X[239:224] * Y[215:192];
            Z53_S1 <= X[223:208] * Y[239:216];
            Z55_S1 <= X[239:224] * Y[239:216];
            Z56_S1 <= X[223:208] * Y[255:240]; // 32 BITS
            Z57_S1 <= X[255:240] * Y[239:216];
            Z58_S1 <= X[239:224] * Y[255:240]; // 32 BITS
            Z60_S1 <= X[255:240] * Y[255:240]; // 32 BITS

            M6_S1 <= (X[15:0] - X[63:48]) * (Y[23:0] - Y[71:48]);
            M8_S1 <= (X[31:16] - X[79:64]) * (Y[23:0] - Y[71:48]);
            M9_S1 <= (X[15:0] - X[63:48]) * (Y[47:24] - Y[95:72]);
            M10_S1 <= (X[47:32] - X[95:80]) * (Y[23:0] - Y[71:48]);
            M11_S1 <= (X[31:16] - X[79:64]) * (Y[47:24] - Y[95:72]);
            M12_S1 <= (X[15:0] - X[111:96]) * (Y[23:0] - Y[119:96]);
            M13_S1 <= (X[47:32] - X[95:80]) * (Y[47:24] - Y[95:72]);
            M14_S1 <= (X[31:16] - X[127:112]) * (Y[23:0] - Y[119:96]);
            M15_S1 <= (X[15:0] - X[111:96]) * (Y[47:24] - Y[143:120]);
            M16_S1 <= (X[47:32] - X[143:128]) * (Y[23:0] - Y[119:96]);
            M17_S1 <= (X[31:16] - X[127:112]) * (Y[47:24] - Y[143:120]);
            M18_0S1 <= (X[63:48] - X[111:96]) * (Y[71:48] - Y[119:96]);
            M18_1S1 <= (X[15:0] - X[159:144]) * (Y[23:0] - Y[167:144]);
            M19_S1 <= (X[47:32] - X[143:128]) * (Y[47:24] - Y[143:120]);
            M20_0S1 <= (X[79:64] - X[127:112]) * (Y[71:48] - Y[119:96]);
            M20_1S1 <= (X[31:16] - X[175:160]) * (Y[23:0] - Y[167:144]);
            M21_0S1 <= (X[15:0] - X[159:144]) * (Y[47:23] - Y[191:168]);
            M21_1S1 <= (X[63:48] - X[111:96]) * (Y[71:48] - Y[119:96]);
            M22_0S1 <= (X[95:80] - X[143:128]) * (Y[71:48] - Y[119:96]);
            M22_1S1 <= (X[47:32] - X[191:176]) * (Y[23:0] - Y[167:144]);
            M23_0S1 <= (X[79:64] - X[127:112]) * (Y[95:72] - Y[143:120]);
            M23_1S1 <= (X[31:16] - X[175:160]) * (Y[47:24] - Y[191:168]);
            M24_0S1 <= (X[15:0] - X[207:192]) * (Y[23:0] - Y[215:192]);
            M24_1S1 <= (X[63:48] - X[159:144]) * (Y[71:48] - Y[167:144]);
            M25_0S1 <= (X[95:80] - X[143:128]) * (Y[95:72] - Y[143:120]);
            M25_1S1 <= (X[47:32] - X[191:176]) * (Y[47:24] - Y[191:168]);
            M26_0S1 <= (X[31:16] - X[223:208]) * (Y[23:0] - Y[215:192]);
            M26_1S1 <= (X[79:64] - X[175:160]) * (Y[71:48] - Y[167:144]);
            M27_0S1 <= (X[15:0] - X[207:192]) * (Y[47:24] - Y[239:216]);
            M27_1S1 <= (X[63:48] - X[159:144]) * (Y[95:72] - Y[191:168]);
            M28_0S1 <= (X[47:32] - X[239:224]) * (Y[23:0] - Y[215:192]);
            M28_1S1 <= (X[95:80] - X[191:176]) * (Y[71:48] - Y[167:144]);
            M29_0S1 <= (X[31:16] - X[223:208]) * (Y[47:24] - Y[239:216]);
            M29_1S1 <= (X[79:64] - X[175:160]) * (Y[95:72] - Y[191:168]);
            M30_0S1 <= (X[15:0] - X[255:240]) * (Y[23:0] - Y[255:240]); 
            M30_1S1 <= (X[63:48] - X[207:192]) * (Y[71:48] - Y[215:192]);
            M30_2S1 <= (X[111:96] - X[159:144]) * (Y[119:96] - Y[167:144]);
            M31_0S1 <= (X[47:32] - X[239:224]) * (Y[47:24] - Y[239:216]);
            M31_1S1 <= (X[95:80] - X[191:176]) * (Y[95:72] - Y[191:168]);
            M32_0S1 <= (X[79:64] - X[175:160]) * (Y[119:96] - Y[215:192]);
            M32_1S1 <= (X[31:16] - X[223:208]) * (Y[71:48] - Y[255:240]);
            M33_0S1 <= (X[63:48] - X[255:240]) * (Y[47:24] - Y[239:216]);
            M33_1S1 <= (X[111:96] - X[207:192]) * (Y[95:72] - Y[191:168]);
            M34_0S1 <= (X[47:32] - X[239:224]) * (Y[71:48] - Y[255:240]);
            M34_1S1 <= (X[95:80] - X[191:176]) * (Y[119:96] - Y[215:192]);
            M35_0S1 <= (X[127:112] - X[175:160]) * (Y[143:120] - Y[191:168]);
            M35_1S1 <= (X[79:64] - X[223:208]) * (Y[95:72] - Y[239:216]);
            M36_0S1 <= (X[63:48] - X[255:240]) * (Y[71:48] - Y[255:240]);
            M36_1S1 <= (X[111:96] - X[207:192]) * (Y[119:96] - Y[215:192]);
            M37_0S1 <= (X[143:128] - X[191:176]) * (Y[143:120] - Y[191:168]);
            M37_1S1 <= (X[95:80] - X[239:224]) * (Y[95:72] - Y[239:216]);
            M38_0S1 <= (X[79:64] - X[223:208]) * (Y[119:96] - Y[255:240]);
            M38_1S1 <= (X[127:112] - X[175:160]) * (Y[167:144] - Y[215:192]);
            M39_0S1 <= (X[111:96] - X[255:240]) * (Y[95:72] - Y[239:216]);
            M39_1S1 <= (X[159:144] - X[207:192]) * (Y[143:120] - Y[191:168]);
            M40_0S1 <= (X[95:80] - X[239:224]) * (Y[119:96] - Y[255:240]);
            M40_1S1 <= (X[143:128] - X[191:176]) * (Y[167:144] - Y[215:192]);
            M41_S1 <= (X[127:112] - X[223:208]) * (Y[143:120] - Y[239:216]);
            M42_0S1 <= (X[159:144] - X[207:192]) * (Y[167:144] - Y[215:192]);
            M42_1S1 <= (X[95:80] - X[239:224]) * (Y[119:96] - Y[255:240]);
            M43_S1 <= (X[143:128] - X[239:224]) * (Y[143:120] - Y[239:216]);
            M44_S1 <= (X[127:112] - X[239:224]) * (Y[167:144] - Y[255:240]);
            M45_S1 <= (X[159:144] - X[255:240]) * (Y[143:120] - Y[239:216]);
            M46_S1 <= (X[143:128] - X[239:224]) * (Y[167:144] - Y[255:240]);
            M47_S1 <= (X[175:160] - X[223:208]) * (Y[191:168] - Y[239:216]);
            M48_S1 <= (X[159:144] - X[255:240]) * (Y[167:144] - Y[255:240]);
            M49_S1 <= (X[191:176] - X[239:224]) * (Y[191:168] - Y[239:216]);
            M50_S1 <= (X[175:160] - X[223:208]) * (Y[215:192] - Y[255:240]);
            M51_S1 <= (X[207:192] - X[255:240]) * (Y[191:168] - Y[239:216]);
            M52_S1 <= (X[191:176] - X[239:224]) * (Y[215:192] - Y[255:240]);
            M54_S1 <= (X[207:192] - X[255:240]) * (Y[215:192] - Y[255:240]);
            
            // Cycle 2
            //S80_0S2 <= Z0_S1 + 


        end
    end

endmodule