`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.08.2025 12:10:40
// Design Name: 
// Module Name: modBRAM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module modBRAM(
    input wire [4:0] type,
    input wire clk,
    input wire start,
    input wire RST,
    output reg [255:0] data,
    output reg done
    );
    
    wire[71:0] DO;
    wire [63:0] DataOut;
    reg[8:0] ADDR;
    reg RDEN;
    
    localparam IDLE = 4'd0, WAIT1 = 4'd1, READ1 = 4'd2, WAIT2 = 4'd3, READ2 = 4'd4, WAIT3 = 4'd5, READ3 = 4'd6, WAIT4 = 4'd7, READ4 = 4'd8, REWAIT1 = 4'd9, REREAD1 = 4'd10;
	assign DataOut = {DO[70:63],DO[61:54],DO[52:45],DO[43:36],DO[34:27],DO[25:18],DO[16:9],DO[7:0]};

    BRAM_SDP_MACRO #(
    .BRAM_SIZE("36Kb"),
    .DEVICE("7SERIES"),
    .WRITE_WIDTH(72),
    .READ_WIDTH(72),
    .DO_REG(0),
    .INIT_FILE("NONE"), // Change to File path before implementation
    .SIM_COLLISION_CHECK("ALL"),
    .SRVAL(72'h00000000000),
    .INIT(72'h00000000000),
    .WRITE_MODE("WRITE_FIRST"),
    
    .INIT_00(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBB),
    .INIT_01(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBB),
    .INIT_02(256'h000000000000000000000),
   .INIT_03(256'h000000000000000000000),
   .INIT_04(256'h000000000000000000000),
   .INIT_05(256'h000000000000000000000),
   .INIT_06(256'h000000000000000000000),
   .INIT_07(256'h000000000000000000000),
   .INIT_08(256'h000000000000000000000),
   .INIT_09(256'h000000000000000000000),
   .INIT_0A(256'h000000000000000000000),
   .INIT_0B(256'h000000000000000000000),
   .INIT_0C(256'h000000000000000000000),
   .INIT_0D(256'h000000000000000000000),
   .INIT_0E(256'h000000000000000000000),
   .INIT_0F(256'h000000000000000000000),
   .INIT_10(256'h000000000000000000000),
   .INIT_11(256'h000000000000000000000),
   .INIT_12(256'h000000000000000000000),
   .INIT_13(256'h000000000000000000000),
   .INIT_14(256'h000000000000000000000),
   .INIT_15(256'h000000000000000000000),
   .INIT_16(256'h000000000000000000000),
   .INIT_17(256'h000000000000000000000),
   .INIT_18(256'h000000000000000000000),
   .INIT_19(256'h000000000000000000000),
   .INIT_1A(256'h000000000000000000000),
   .INIT_1B(256'h000000000000000000000),
   .INIT_1C(256'h000000000000000000000),
   .INIT_1D(256'h000000000000000000000),
   .INIT_1E(256'h000000000000000000000),
   .INIT_1F(256'h000000000000000000000),
   .INIT_20(256'h000000000000000000000),
   .INIT_21(256'h000000000000000000000),
   .INIT_22(256'h000000000000000000000),
   .INIT_23(256'h000000000000000000000),
   .INIT_24(256'h000000000000000000000),
   .INIT_25(256'h000000000000000000000),
   .INIT_26(256'h000000000000000000000),
   .INIT_27(256'h000000000000000000000),
   .INIT_28(256'h000000000000000000000),
   .INIT_29(256'h000000000000000000000),
   .INIT_2A(256'h000000000000000000000),
   .INIT_2B(256'h000000000000000000000),
   .INIT_2C(256'h000000000000000000000),
   .INIT_2D(256'h000000000000000000000),
   .INIT_2E(256'h000000000000000000000),
   .INIT_2F(256'h000000000000000000000),
   .INIT_30(256'h000000000000000000000),
   .INIT_31(256'h000000000000000000000),
   .INIT_32(256'h000000000000000000000),
   .INIT_33(256'h000000000000000000000),
   .INIT_34(256'h000000000000000000000),
   .INIT_35(256'h000000000000000000000),
   .INIT_36(256'h000000000000000000000),
   .INIT_37(256'h000000000000000000000),
   .INIT_38(256'h000000000000000000000),
   .INIT_39(256'h000000000000000000000),
   .INIT_3A(256'h000000000000000000000),
   .INIT_3B(256'h000000000000000000000),
   .INIT_3C(256'h000000000000000000000),
   .INIT_3D(256'h000000000000000000000),
   .INIT_3E(256'h000000000000000000000),
   .INIT_3F(256'h000000000000000000000),

   // The next set of INIT_xx are valid when configured as 36Kb
   .INIT_40(256'h000000000000000000000),
   .INIT_41(256'h000000000000000000000),
   .INIT_42(256'h000000000000000000000),
   .INIT_43(256'h000000000000000000000),
   .INIT_44(256'h000000000000000000000),
   .INIT_45(256'h000000000000000000000),
   .INIT_46(256'h000000000000000000000),
   .INIT_47(256'h000000000000000000000),
   .INIT_48(256'h000000000000000000000),
   .INIT_49(256'h000000000000000000000),
   .INIT_4A(256'h000000000000000000000),
   .INIT_4B(256'h000000000000000000000),
   .INIT_4C(256'h000000000000000000000),
   .INIT_4D(256'h000000000000000000000),
   .INIT_4E(256'h000000000000000000000),
   .INIT_4F(256'h000000000000000000000),
   .INIT_50(256'h000000000000000000000),
   .INIT_51(256'h000000000000000000000),
   .INIT_52(256'h000000000000000000000),
   .INIT_53(256'h000000000000000000000),
   .INIT_54(256'h000000000000000000000),
   .INIT_55(256'h000000000000000000000),
   .INIT_56(256'h000000000000000000000),
   .INIT_57(256'h000000000000000000000),
   .INIT_58(256'h000000000000000000000),
   .INIT_59(256'h000000000000000000000),
   .INIT_5A(256'h000000000000000000000),
   .INIT_5B(256'h000000000000000000000),
   .INIT_5C(256'h000000000000000000000),
   .INIT_5D(256'h000000000000000000000),
   .INIT_5E(256'h000000000000000000000),
   .INIT_5F(256'h000000000000000000000),
   .INIT_60(256'h000000000000000000000),
   .INIT_61(256'h000000000000000000000),
   .INIT_62(256'h000000000000000000000),
   .INIT_63(256'h000000000000000000000),
   .INIT_64(256'h000000000000000000000),
   .INIT_65(256'h000000000000000000000),
   .INIT_66(256'h000000000000000000000),
   .INIT_67(256'h000000000000000000000),
   .INIT_68(256'h000000000000000000000),
   .INIT_69(256'h000000000000000000000),
   .INIT_6A(256'h000000000000000000000),
   .INIT_6B(256'h000000000000000000000),
   .INIT_6C(256'h000000000000000000000),
   .INIT_6D(256'h000000000000000000000),
   .INIT_6E(256'h000000000000000000000),
   .INIT_6F(256'h000000000000000000000),
   .INIT_70(256'h000000000000000000000),
   .INIT_71(256'h000000000000000000000),
   .INIT_72(256'h000000000000000000000),
   .INIT_73(256'h000000000000000000000),
   .INIT_74(256'h000000000000000000000),
   .INIT_75(256'h000000000000000000000),
   .INIT_76(256'h000000000000000000000),
   .INIT_77(256'h000000000000000000000),
   .INIT_78(256'h000000000000000000000),
   .INIT_79(256'h000000000000000000000),
   .INIT_7A(256'h000000000000000000000),
   .INIT_7B(256'h000000000000000000000),
   .INIT_7C(256'h000000000000000000000),
   .INIT_7D(256'h000000000000000000000),
   .INIT_7E(256'h000000000000000000000),
   .INIT_7F(256'h000000000000000000000),

   // The next set of INITP_xx are for the parity bits
   .INITP_00(256'h000000000000000000000),
   .INITP_01(256'h000000000000000000000),
   .INITP_02(256'h000000000000000000000),
   .INITP_03(256'h000000000000000000000),
   .INITP_04(256'h000000000000000000000),
   .INITP_05(256'h000000000000000000000),
   .INITP_06(256'h000000000000000000000),
   .INITP_07(256'h000000000000000000000),

   // The next set of INITP_xx are valid when configured as 36Kb
   .INITP_08(256'h000000000000000000000),
   .INITP_09(256'h000000000000000000000),
   .INITP_0A(256'h000000000000000000000),
   .INITP_0B(256'h000000000000000000000),
   .INITP_0C(256'h000000000000000000000),
   .INITP_0D(256'h000000000000000000000),
   .INITP_0E(256'h000000000000000000000),
   .INITP_0F(256'h000000000000000000000) 
    ) BRAM_SDP_MACRO_inst (
    .DO(DO),
    .DI(72'h00000000000000000),
    .RDADDR(ADDR),
    .RDCLK(clk),
    .RDEN(RDEN),
    .REGCE(1'b1),
    .RST(RST),
    .WE(8'h00),
    .WRADDR(ADDR),
    .WRCLK(clk),
    .WREN(0)
    );
    
    reg [3:0] state;
    
    always @(posedge clk) begin
    	if(RST) begin
    		done <= 0;
    		RDEN <= 0;
    		data <= 0;
    		state <= IDLE;
    		ADDR <= 9'b110000000;
		end  		
    	
		case(state) 
			IDLE: begin
				done <= 0;
				RDEN <= 0;
				if(start) begin
					state <= WAIT1;
					RDEN <= 1;
					ADDR <= {2'b00, type, 2'b00};
				end
			end
			
			WAIT1: begin
				state <= READ1;
				RDEN <= 0;
			end
			
			READ1: begin
				ADDR <= {2'b00, type, 2'b01};
				data[63:0] <= DataOut;
				RDEN <= 1;
				state <= WAIT2;
			end
			
			WAIT2: begin
				state <= READ2;
				RDEN <= 0;
			end
			
			READ2: begin
				ADDR <= {2'b00, type, 2'b10};
				RDEN <= 1;
				data[127:64] <= DataOut;
				state <= WAIT3;
			end
			
			WAIT3: begin	
				state <= READ3;
				RDEN <= 0;
			end
			
			READ3: begin
				ADDR <= {2'b00, type, 2'b11};
				data[191:128] <= DataOut;
				RDEN <= 1;
				state <= WAIT4;
			end
			
			WAIT4: begin
				RDEN <= 0;
				state <= READ4;
			end
			
			READ4: begin
				ADDR <= {2'b00, type, 2'b00};
				data[255:192] <= DataOut;
				RDEN <= 1;
				state <= REWAIT1;
			end
			
			REWAIT1: begin
				RDEN <= 0;
				state <= REREAD1;
			end
			
			REREAD1: begin
				data[63:0] <= DataOut;
				done <= 1;
				state <= IDLE;
			end
			
			default: state <= IDLE;
		endcase
	end    			
endmodule 