`timescale 1ns/1ps

module fastKaratsuba(
    input wire clock,
    input wire reset,
    input wire [255:0] X,
    input wire [255:0] Y,
    input wire in_valid,
    output reg [511:0] P,
    output reg out_valid
);

    // Cycle 1
    reg [39:0] Z0_S1, Z2_S1, Z3_S1, Z4_S1, Z5_S1, Z7_S1, Z8_S1, Z9_S1,
                Z10_S1, Z12_S1, Z14_S1, Z15_S1, Z16_S1, Z17_S1, Z19_S1,
                Z20_S1, Z21_S1, Z22_S1, Z24_S1, Z26_S1, Z27_S1, Z28_S1, Z29_S1,
                Z31_S1, Z32_S1, Z33_S1, Z34_S1, Z36_S1, Z38_S1, Z39_S1,
                Z40_S1, Z41_S1, Z43_S1, Z44_S1, Z45_S1, Z46_S1, Z48_S1,
                Z50_S1, Z51_S1, Z52_S1, Z53_S1, Z55_S1, Z57_S1;
    reg [31:0] Z56_S1, Z58_S1, Z60_S1;

    reg [40:0] M6_S1, M8_S1, M9_S1, M10_S1, M11_S1, M12_S1, M13_S1, M14_S1, M15_S1, M16_S1, M17_S1, M18_0S1, M18_1S1, M19_S1,
                M20_0S1, M20_1S1, M21_0S1, M21_1S1, M22_0S1, M22_1S1, M23_0S1, M23_1S1, M24_0S1, M24_1S1, M25_0S1, M25_1S1,
                M26_0S1, M26_1S1, M27_0S1, M27_1S1, M28_0S1, M28_1S1, M29_0S1, M29_1S1, M30_0S1, M30_1S1, M30_2S1, M31_0S1,
                M31_1S1, M32_0S1, M32_1S1, M33_0S1, M33_1S1, M34_0S1, M34_1S1, M35_0S1, M35_1S1, M36_0S1, M36_1S1, M37_0S1,
                M37_1S1, M38_0S1, M38_1S1, M39_0S1, M39_1S1, M40_0S1, M40_1S1, M41_S1, M42_0S1, M42_1S1, M43_S1, M44_S1, M45_S1,
                M46_S1, M47_S1, M48_S1, M49_S1, M50_S1, M51_S1, M52_S1, M54_S1; 
    reg S1_valid;

    // Cycle 2
    reg [80:0] S80_0S2;
    reg [57:0] S106_48S2;
    reg [56:0] S489_432S2; 
    reg [54:0] S511_456S2;
    reg [50:0] S139_88S2, S155_104S2, S171_120S2, S195_144S2, S387_336S2, S403_352S2, S465_416S2;
    reg [49:0] S122_72S2, S186_136S2, S378_328S2, S418_368S2, S434_384S2, S450_400S2;
    reg [42:0] S203_160S2, S211_168S2, S219_176S2, S227_184S2, S235_192S2, S243_200S2, S251_208S2, S259_216S2, S267_224S2, S275_232S2, S283_240S2,
                S291_248S2, S299_256S2, S307_264S2, S315_272S2, S323_280S2, S331_288S2, S339_296S2, S347_304S2, S355_312S2, S363_320S2;

    reg S2_valid;

    // Cycle 3
    reg [123:0] S123_0S3;
    reg [98:0] S187_88S3, S451_352S3;
    reg [94:0] S511_416S3;
    reg [75:0] S220_144S3, S388_312S3;
    reg [67:0] S252_184S3, S284_216S3, S316_248S3, S348_280S3;
    
    reg S3_valid;

    // Cycle 4
    reg [188:0] S188_0S4;
    reg [158:0] S511_352S4;
    reg [108:0] S253_144S4, S389_280S4;
    reg [100:0] S317_216S4;

    reg S4_valid;

    // Cycle 5
    reg [254:0] S254_0S5;
    reg [173:0] S390_216S5;
    reg [158:0] S511_352S5;

    reg S5_valid;

    // Cycle 6
    reg [391:0] S391_0S6;
    reg [158:0] S511_352S6;

    reg S6_valid;

    always @(posedge clock) begin
        if(reset) begin
            P <= 256'b0;
            S1_valid <= 1'b0;
            S2_valid <= 1'b0;
            S3_valid <= 1'b0;
            out_valid <= 1'b0;
        end
        else begin

            // Cycle 1
            Z0_S1 <= X[15:0] * Y[23:0];
            Z2_S1 <= X[31:16] * Y[23:0];
            Z3_S1 <= X[15:0] * Y[47:24];
            Z4_S1 <= X[47:32] * Y[23:0];
            Z5_S1 <= X[31:16] * Y[47:24];
            Z7_S1 <= X[47:32] * Y[47:24];
            Z8_S1 <= X[31:16] * Y[71:48];
            Z9_S1 <= X[63:48] * Y[47:24];
            Z10_S1 <= X[47:32] * Y[71:48];
            Z12_S1 <= X[63:48] * Y[71:48];
            Z14_S1 <= X[79:64] * Y[71:48];
            Z15_S1 <= X[63:48] * Y[95:72];
            Z16_S1 <= X[97:80] * Y[71:48];
            Z17_S1 <= X[79:64] * Y[95:72];
            Z19_S1 <= X[95:80] * Y[95:72];
            Z20_S1 <= X[79:64] * Y[119:96];
            Z21_S1 <= X[111:96] * Y[95:72];
            Z22_S1 <= X[95:80] * Y[119:96];
            Z24_S1 <= X[111:96] * Y[119:96];
            Z26_S1 <= X[127:112] * Y[119:96];
            Z27_S1 <= X[111:96] * Y[143:120];
            Z28_S1 <= X[143:128] * Y[119:96];
            Z29_S1 <= X[127:112] * Y[143:120];
            Z31_S1 <= X[143:128] * Y[143:120];
            Z32_S1 <= X[127:112] * Y[167:144];
            Z33_S1 <= X[159:144] * Y[143:120];
            Z34_S1 <= X[143:128] * Y[167:144];
            Z36_S1 <= X[159:144] * Y[167:144];
            Z38_S1 <= X[175:160] * Y[167:144];
            Z39_S1 <= X[159:144] * Y[191:168];
            Z40_S1 <= X[191:176] * Y[167:144];
            Z41_S1 <= X[175:160] * Y[191:168];
            Z43_S1 <= X[191:176] * Y[191:168];
            Z44_S1 <= X[175:160] * Y[215:192];
            Z45_S1 <= X[207:192] * Y[191:168];
            Z46_S1 <= X[191:176] * Y[215:192];
            Z48_S1 <= X[207:192] * Y[215:192];
            Z50_S1 <= X[223:208] * Y[215:192];
            Z51_S1 <= X[207:192] * Y[239:216];
            Z52_S1 <= X[239:224] * Y[215:192];
            Z53_S1 <= X[223:208] * Y[239:216];
            Z55_S1 <= X[239:224] * Y[239:216];
            Z56_S1 <= X[223:208] * Y[255:240]; // 32 BITS
            Z57_S1 <= X[255:240] * Y[239:216];
            Z58_S1 <= X[239:224] * Y[255:240]; // 32 BITS
            Z60_S1 <= X[255:240] * Y[255:240]; // 32 BITS

            M6_S1 <= ($signed({1'b0, X[15:0]}) - $signed({1'b0, X[63:48]})) * ($signed({1'b0, Y[71:48]}) - $signed({1'b0, Y[23:0]}));
            M8_S1 <= (X[31:16] - X[79:64]) * ( - Y[23:0] + Y[71:48]);
            M9_S1 <= (X[15:0] - X[63:48]) * ( - Y[47:24] + Y[95:72]);
            M10_S1 <= (X[47:32] - X[95:80]) * ( - Y[23:0] + Y[71:48]);
            M11_S1 <= (X[31:16] - X[79:64]) * ( - Y[47:24] + Y[95:72]);
            M12_S1 <= (X[15:0] - X[111:96]) * ( - Y[23:0] + Y[119:96]);
            M13_S1 <= (X[47:32] - X[95:80]) * ( - Y[47:24] + Y[95:72]);
            M14_S1 <= (X[31:16] - X[127:112]) * ( - Y[23:0] + Y[119:96]);
            M15_S1 <= (X[15:0] - X[111:96]) * ( - Y[47:24] + Y[143:120]);
            M16_S1 <= (X[47:32] - X[143:128]) * ( - Y[23:0] + Y[119:96]);
            M17_S1 <= (X[31:16] - X[127:112]) * ( - Y[47:24] + Y[143:120]);
            M18_0S1 <= (X[63:48] - X[111:96]) * ( - Y[71:48] + Y[119:96]);
            M18_1S1 <= (X[15:0] - X[159:144]) * ( - Y[23:0] + Y[167:144]);
            M19_S1 <= (X[47:32] - X[143:128]) * ( - Y[47:24] + Y[143:120]);
            M20_0S1 <= (X[79:64] - X[127:112]) * ( - Y[71:48] + Y[119:96]);
            M20_1S1 <= (X[31:16] - X[175:160]) * ( - Y[23:0] + Y[167:144]);
            M21_0S1 <= (X[15:0] - X[159:144]) * ( - Y[47:23] + Y[191:168]);
            M21_1S1 <= (X[63:48] - X[111:96]) * ( - Y[71:48] + Y[119:96]);
            M22_0S1 <= (X[95:80] - X[143:128]) * ( - Y[71:48] + Y[119:96]);
            M22_1S1 <= (X[47:32] - X[191:176]) * ( - Y[23:0] + Y[167:144]);
            M23_0S1 <= (X[79:64] - X[127:112]) * ( - Y[95:72] + Y[143:120]);
            M23_1S1 <= (X[31:16] - X[175:160]) * ( - Y[47:24] + Y[191:168]);
            M24_0S1 <= (X[15:0] - X[207:192]) * ( - Y[23:0] + Y[215:192]);
            M24_1S1 <= (X[63:48] - X[159:144]) * ( - Y[71:48] + Y[167:144]);
            M25_0S1 <= (X[95:80] - X[143:128]) * ( - Y[95:72] + Y[143:120]);
            M25_1S1 <= (X[47:32] - X[191:176]) * ( - Y[47:24] + Y[191:168]);
            M26_0S1 <= (X[31:16] - X[223:208]) * ( - Y[23:0] + Y[215:192]);
            M26_1S1 <= (X[79:64] - X[175:160]) * ( - Y[71:48] + Y[167:144]);
            M27_0S1 <= (X[15:0] - X[207:192]) * ( - Y[47:24] + Y[239:216]);
            M27_1S1 <= (X[63:48] - X[159:144]) * ( - Y[95:72] + Y[191:168]);
            M28_0S1 <= (X[47:32] - X[239:224]) * ( - Y[23:0] + Y[215:192]);
            M28_1S1 <= (X[95:80] - X[191:176]) * ( - Y[71:48] + Y[167:144]);
            M29_0S1 <= (X[31:16] - X[223:208]) * ( - Y[47:24] + Y[239:216]);
            M29_1S1 <= (X[79:64] - X[175:160]) * ( - Y[95:72] + Y[191:168]);
            M30_0S1 <= (X[15:0] - X[255:240]) * ( - Y[23:0] + Y[255:240]); 
            M30_1S1 <= (X[63:48] - X[207:192]) * ( - Y[71:48] + Y[215:192]);
            M30_2S1 <= (X[111:96] - X[159:144]) * ( - Y[119:96] + Y[167:144]);
            M31_0S1 <= (X[47:32] - X[239:224]) * ( - Y[47:24] + Y[239:216]);
            M31_1S1 <= (X[95:80] - X[191:176]) * ( - Y[95:72] + Y[191:168]);
            M32_0S1 <= (X[79:64] - X[175:160]) * ( - Y[119:96] + Y[215:192]);
            M32_1S1 <= (X[31:16] - X[223:208]) * ( - Y[71:48] + Y[255:240]);
            M33_0S1 <= (X[63:48] - X[255:240]) * ( - Y[47:24] + Y[239:216]);
            M33_1S1 <= (X[111:96] - X[207:192]) * ( - Y[95:72] + Y[191:168]);
            M34_0S1 <= (X[47:32] - X[239:224]) * ( - Y[71:48] + Y[255:240]);
            M34_1S1 <= (X[95:80] - X[191:176]) * ( - Y[119:96] + Y[215:192]);
            M35_0S1 <= (X[127:112] - X[175:160]) * ( - Y[143:120] + Y[191:168]);
            M35_1S1 <= (X[79:64] - X[223:208]) * ( - Y[95:72] + Y[239:216]);
            M36_0S1 <= (X[63:48] - X[255:240]) * ( - Y[71:48] + Y[255:240]);
            M36_1S1 <= (X[111:96] - X[207:192]) * ( - Y[119:96] + Y[215:192]);
            M37_0S1 <= (X[143:128] - X[191:176]) * ( - Y[143:120] + Y[191:168]);
            M37_1S1 <= (X[95:80] - X[239:224]) * ( - Y[95:72] + Y[239:216]);
            M38_0S1 <= (X[79:64] - X[223:208]) * ( - Y[119:96] + Y[255:240]);
            M38_1S1 <= (X[127:112] - X[175:160]) * ( - Y[167:144] + Y[215:192]);
            M39_0S1 <= (X[111:96] - X[255:240]) * ( - Y[95:72] + Y[239:216]);
            M39_1S1 <= (X[159:144] - X[207:192]) * ( - Y[143:120] + Y[191:168]);
            M40_0S1 <= (X[95:80] - X[239:224]) * ( - Y[119:96] + Y[255:240]);
            M40_1S1 <= (X[143:128] - X[191:176]) * ( - Y[167:144] + Y[215:192]);
            M41_S1 <= (X[127:112] - X[223:208]) * ( - Y[143:120] + Y[239:216]);
            M42_0S1 <= (X[159:144] - X[207:192]) * ( - Y[167:144] + Y[215:192]);
            M42_1S1 <= (X[95:80] - X[239:224]) * ( - Y[119:96] + Y[255:240]);
            M43_S1 <= (X[143:128] - X[239:224]) * ( - Y[143:120] + Y[239:216]);
            M44_S1 <= (X[127:112] - X[239:224]) * ( - Y[167:144] + Y[255:240]);
            M45_S1 <= (X[159:144] - X[255:240]) * ( - Y[143:120] + Y[239:216]);
            M46_S1 <= (X[143:128] - X[239:224]) * ( - Y[167:144] + Y[255:240]);
            M47_S1 <= (X[175:160] - X[223:208]) * ( - Y[191:168] + Y[239:216]);
            M48_S1 <= (X[159:144] - X[255:240]) * ( - Y[167:144] + Y[255:240]);
            M49_S1 <= (X[191:176] - X[239:224]) * ( - Y[191:168] + Y[239:216]);
            M50_S1 <= (X[175:160] - X[223:208]) * ( - Y[215:192] + Y[255:240]);
            M51_S1 <= (X[207:192] - X[255:240]) * ( - Y[191:168] + Y[239:216]);
            M52_S1 <= (X[191:176] - X[239:224]) * ( - Y[215:192] + Y[255:240]);
            M54_S1 <= (X[207:192] - X[255:240]) * ( - Y[215:192] + Y[255:240]);
            
            S1_valid <= in_valid;
            
            // Cycle 2
            S80_0S2 <= Z0_S1 + {Z2_S1, 16'b0} + {Z3_S1, 24'b0} + {Z4_S1, 32'b0} + {Z5_S1, 40'b1};
            S106_48S2 <= M6_S1 + Z0_S1 + Z12_S1 + {Z7_S1, 8'b0} + {M8_S1, 16'b0} + {Z2_S1, 16'b0} + {Z14_S1, 16'b0};
            S122_72S2 <= M9_S1 + Z3_S1 + Z15_S1 + {M10_S1, 8'b0} + {Z4_S1, 8'b0} + {Z16_S1, 8'b0};
            S139_88S2 <= M11_S1 + Z5_S1 + Z17_S1 + {Z12_S1, 8'b0} + {M12_S1, 8'b0} + {Z0_S1, 8'b0} + {Z24_S1, 8'b0};
            S155_104S2 <= M13_S1 + Z7_S1 + Z19_S1 + {Z14_S1, 8'b0} + {M14_S1, 8'b0} + {Z2_S1, 8'b0} + {Z26_S1, 8'b0};
            S171_120S2 <= Z15_S1 + M15_S1 + Z3_S1 + Z27_S1 + {Z16_S1, 8'b0} + {M16_S1, 8'b0} + {Z4_S1, 8'b0} + {Z28_S1, 8'b0};
            S186_136S2 <= Z17_S1 + M17_S1 + Z5_S1 + Z29_S1 + {M18_0S1, 8'b0} + {Z12_S1, 8'b0} + {Z24_S1, 8'b0};
            S195_144S2 <= M18_1S1 + Z0_S1 + Z36_S1 + {Z19_S1, 8'b0} + {M19_S1, 8'b0} + {Z7_S1, 8'b0} + {Z31_S1, 8'b0};
            S203_160S2 <= M20_0S1 + M20_1S1 + Z14_S1 + Z26_S1 + Z2_S1 + Z38_S1;
            S211_168S2 <= M21_0S1 + M21_1S1 + Z15_S1 + Z27_S1 + Z3_S1 + Z39_S1;
            S219_176S2 <= M22_0S1 + M22_1S1 + Z16_S1 + Z28_S1 + Z4_S1 + Z40_S1;
            S227_184S2 <= M23_0S1 + M23_1S1 + Z17_S1 + Z29_S1 + Z5_S1 + Z41_S1;
            S235_192S2 <= M24_0S1 + M24_1S1 + Z24_S1 + Z12_S1 + Z36_S1 + Z0_S1 + Z48_S1;
            S243_200S2 <= M25_0S1 + M25_1S1 + Z19_S1 + Z31_S1 + Z7_S1 + Z43_S1;
            S251_208S2 <= M26_0S1 + M26_1S1 + Z26_S1 + Z14_S1 + Z38_S1 + Z2_S1 + Z50_S1;
            S259_216S2 <= M27_0S1 + M27_1S1 + Z27_S1 + Z15_S1 + Z39_S1 + Z3_S1 + Z51_S1;
            S267_224S2 <= M28_0S1 + M28_1S1 + Z28_S1 + Z16_S1 + Z40_S1 + Z4_S1 + Z52_S1;
            S275_232S2 <= M29_0S1 + M29_1S1 + Z29_S1 + Z17_S1 + Z41_S1 + Z5_S1 + Z53_S1;
            S283_240S2 <= M30_0S1 + M30_1S1 + M30_2S1 + Z0_S1 + Z12_S1 + Z24_S1 + Z36_S1 + Z48_S1 + Z60_S1;
            S291_248S2 <= M31_0S1 + M31_1S1 + Z31_S1 + Z19_S1 + Z43_S1 + Z7_S1 + Z55_S1;
            S299_256S2 <= M32_0S1 + M32_1S1 + Z32_S1 + Z20_S1 + Z44_S1 + Z8_S1 + Z56_S1;
            S307_264S2 <= M33_0S1 + M33_1S1 + Z33_S1 + Z21_S1 + Z45_S1 + Z9_S1 + Z57_S1;
            S315_272S2 <= M34_0S1 + M34_1S1 + Z34_S1 + Z22_S1 + Z46_S1 + Z10_S1 + Z58_S1;
            S323_280S2 <= M35_0S1 + M35_1S1 + Z29_S1 + Z41_S1 + Z17_S1 + Z53_S1;
            S331_288S2 <= M36_0S1 + M36_1S1 + Z36_S1 + Z12_S1 + Z24_S1 + Z48_S1 + Z60_S1;
            S339_296S2 <= M37_0S1 + M37_1S1 + Z31_S1 + Z43_S1 + Z19_S1 + Z55_S1;
            S347_304S2 <= M38_0S1 + M38_1S1 + Z32_S1 + Z44_S1 + Z20_S1 + Z56_S1;
            S355_312S2 <= M39_0S1 + M39_1S1 + Z33_S1 + Z45_S1 + Z21_S1 + Z57_S1;
            S363_320S2 <= M40_0S1 + M40_1S1 + Z34_S1 + Z46_S1 + Z22_S1 + Z58_S1;
            S378_328S2 <= M41_S1 + Z41_S1 + Z29_S1 + Z53_S1 + {M42_0S1, 8'b0} + {Z36_S1, 8'b0} + {Z48_S1, 8'b0};
            S387_336S2 <= M42_1S1 + Z24_S1 + Z60_S1 + {M43_S1, 8'b0} + {Z43_S1, 8'b0} + {Z31_S1, 8'b0} + {Z53_S1, 8'b0};
            S403_352S2 <= M44_S1 + Z44_S1 + Z32_S1 + Z56_S1 + {M45_S1, 8'b0} + {Z45_S1, 8'b0} + {Z33_S1, 8'b0} + {Z57_S1, 8'b0};
            S418_368S2 <= M46_S1 + Z46_S1 + Z34_S1 + Z58_S1 + {M47_S1, 8'b0} + {Z41_S1, 8'b0} + {Z53_S1, 8'b0};
            S434_384S2 <= M48_S1 + Z48_S1 + Z36_S1 + Z60_S1 + {M49_S1, 8'b0} + {Z43_S1, 8'b0} + {Z55_S1, 8'b0};
            S450_400S2 <= M50_S1 + Z44_S1 + Z56_S1 + {M51_S1, 8'b0} + {Z45_S1, 8'b0} + {Z57_S1, 8'b0};
            S465_416S2 <= M52_S1 + Z46_S1 + Z58_S1 + {Z53_S1, 8'b0};
            S489_432S2 <= M54_S1 + Z48_S1 + Z60_S1 + {Z55_S1, 8'b0} + {Z56_S1, 16'b0};
            S511_456S2 <= Z57_S1 + {Z58_S1, 8'b0} + {Z60_S1, 24'b0};

            S2_valid <= S1_valid;

            // Cycle 3
            S123_0S3 <= S80_0S2 + {S106_48S2, 48'b0} + {S122_72S2, 72'b0};
            S187_88S3 <= S139_88S2 + {S155_104S2, 16'b0} + {S171_120S2, 32'b0} + {S186_136S2, 48'b0};
            S220_144S3 <= S195_144S2 + {S203_160S2, 16'b0} + {S211_168S2, 24'b0} + {S219_176S2, 32'b0};
            S252_184S3 <= S227_184S2 + {S235_192S2, 8'b0} + {S243_200S2, 16'b0} + {S251_208S2, 24'b0};
            S284_216S3 <= S259_216S2 + {S267_224S2, 8'b0} + {S275_232S2, 16'b0} + {S283_240S2, 24'b0};
            S316_248S3 <= S291_248S2 + {S299_256S2, 8'b0} + {S307_264S2, 16'b0} + {S315_272S2, 24'b0};
            S348_280S3 <= S323_280S2 + {S331_288S2, 8'b0} + {S339_296S2, 16'b0} + {S347_304S2, 24'b0};
            S388_312S3 <= S355_312S2 + {S363_320S2, 8'b0} + {S378_328S2, 16'b0} + {S387_336S2, 24'b0};
            S451_352S3 <= S403_352S2 + {S418_368S2, 16'b0} + {S434_384S2, 32'b0} + {S450_400S2, 48'b0};
            S511_416S3 <= S465_416S2 + {S489_432S2, 16'b0} + {S511_456S2, 40'b0};

            S3_valid <= S2_valid;

            // Cycle 4 
            S188_0S4 <= S123_0S3 + {S187_88S3, 88'b0};
            S253_144S4 <= S220_144S3 + {S252_184S3, 40'b0};
            S317_216S4 <= S284_216S3 + {S316_248S3, 32'b0};
            S389_280S4 <= S348_280S3 + {S388_312S3, 32'b0};
            S511_352S4 <= S451_352S3 + {S511_416S3, 64'b0};

            S4_valid <= S3_valid;

            // Cycle 5
            S254_0S5 <= S188_0S4 + {S253_144S4, 144'b0};
            S390_216S5 <= S317_216S4 + {S389_280S4, 64'b0};
            S511_352S5 <= S511_352S4;

            S5_valid <= S4_valid;

            // Cycle 6
            S391_0S6 <= S254_0S5 + {S390_216S5, 216'b0};
            S511_352S6 <= S511_352S5;

            S6_valid <= S5_valid;

            // Cycle 7
            P <= S391_0S6 + {S511_352S6, 352'b0};

            out_valid <= S6_valid;
        end
    end

endmodule